

 
 
 




window new WaveWindow  -name  "Waves for BMG Example Design"
waveform  using  "Waves for BMG Example Design"

      waveform add -signals /I_RAM_tb/status
      waveform add -signals /I_RAM_tb/I_RAM_synth_inst/bmg_port/CLKA
      waveform add -signals /I_RAM_tb/I_RAM_synth_inst/bmg_port/ADDRA
      waveform add -signals /I_RAM_tb/I_RAM_synth_inst/bmg_port/DINA
      waveform add -signals /I_RAM_tb/I_RAM_synth_inst/bmg_port/WEA
      waveform add -signals /I_RAM_tb/I_RAM_synth_inst/bmg_port/DOUTA

console submit -using simulator -wait no "run"
